///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: MUX2_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"

///////////////////////////////////////////////////////////////////////////////////
// Inputs: A, B (32-bit); S (1-bit)
reg[31:0] A;
reg[31:0] B;
reg S;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Output: Y (32-bit)
wire[31:0] Y;
///////////////////////////////////////////////////////////////////////////////////

MUX2_32 myMUX(.S(S), 
              .A(A), 
              .B(B), 
              .Y(Y));

initial begin
/////////////////////////////////////////////////////////////////////////////
// Test: S=0
$display("Testing S=0: ");
A=32767; B=25879; S=0;  #10; 
verifyEqual32(Y, A);
/////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////
// Test: S=1
$display("Testing S=1: ");
S=1;  #10; 
verifyEqual32(Y, B);
/////////////////////////////////////////////////////////////////////////////
$display("All tests passed.");
end

endmodule